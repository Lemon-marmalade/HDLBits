module top_module(
    input clk,
    input load,
    input [255:0] data,
    output [255:0] q ); 
    
    reg [255:0] q_next;
    integer i, j;
    integer i_s, i_a, j_s, j_a;
    // this solution is a bit manual and tedious, fix this some time
    always @(*) begin
        for(i = 0; i < 16; ++ i)
            for(j = 0; j < 16; ++ j)
                begin
                    if(i == 0)
                        i_s = 15; // right of right edge
                    else
                        i_s = i - 1;
                    
                    if(j == 0)
                        j_s = 15; //bottom of bottom edge
                    else
                        j_s = j - 1;
                    
                    if(i == 15)
                        i_a = 0; // left of left edge
                    else
                        i_a = i + 1;
                    
                    if(j == 15)
                        j_a = 0; // top of top edge
                    else
                        j_a = j + 1;
                    
                    case(q[i_a+j_s*16] + q[i_s+j_a*16] + q[i_s+j_s*16] + q[i_a+j_a*16] + q[i_s+j*16] + q[i_a+j*16] + q[i+j_s*16] + q[i+j_a*16])
                        4'b0010: q_next[i+j*16] <= q[i+j*16];
                        4'b0011: q_next[i+j*16] <= 1;
                        default: q_next[i+j*16] <= 0;
                    endcase
                end
    end
    
    always @(posedge clk) begin
        if(load)
            q <= data;
        else
	    	q <= q_next;
    end

endmodule

/* Revisiting Conway's Game of Life (to fix very delicate and unstable edge case logic from before)

module top_module(
    input clk,
    input load,
    input [255:0] data,
    output [255:0] q ); 
    
    integer i, j;
    integer l, r, t, b, n;
    reg [255:0] next_q;
    
    always @(*) begin
        for (i=0;i<16;i++) begin
            for (j=0; j<16;j++) begin
                // Precalculate edge cases
                l= (j==0)? 15:(j-1);
                r = (j==15)? 0:(j+1);
                b = (i==0)? 15:(i-1);
                t = (i==15)? 0:(i+1);
                // Calculate how many neighbours
                n = (q[i*16+l]+q[t*16+l]+q[t*16+j]+q[t*16+r]+q[i*16+r]+q[b*16+r]+q[b*16+j]+q[b*16+l]);

                if (n<2||n>3)
                    next_q[i*16+j]<=0;
                else if (n==3)
                    next_q[i*16+j]<=1;
                else
                    next_q[i*16+j]<=q[i*16+j];
            end
        end
    end
    
    always @(posedge clk) begin
        if (load)
            q<=data;
        else
            q<=next_q;
    end
    
endmodule

*/
