module top_module (
    input clk,
    input reset,        // Synchronous active-high reset
    output [3:0] q);
    
    always @ (posedge clk) begin
        if (reset || q==9)
            q <= 4'b0;
        else
            q <= q + 4'h1;
    end

endmodule